`define OP_NULL    3'h0
`define OP_ADD     3'h1
`define OP_SUB     3'h2
`define OP_MUL     3'h3
`define OP_DIV     3'h4
`define OP_AND     3'h5
`define OP_LEFT3   3'h6
`define OP_LEFT4   3'h7